// 
// ${copyright_header}
// Copyright 2020 Datum Technology Corporation
// 
// Licensed under the Solderpad Hardware License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
// 
//     https://solderpad.org/licenses/
// 
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// 


`ifndef __UVME_${name_uppercase}_CHKR_SV__
`define __UVME_${name_uppercase}_CHKR_SV__


/**
 * TODO Describe uvme_${name}_chkr
 */
module uvme_${name}_chkr (
   // TODO Add interfaces to uvme_${name}_chkr
);
   
   `pragma protect begin
   
   // TODO Add assertions to uvma_reset_if_chkr
   
   `pragma protect end
   
endmodule : uvme_${name}_chkr


`endif // __UVME_${name_uppercase}_CHKR_SV__
